module reorder_buffer(
	//inputs: 2 inputs; 1 from address unit, 1 from CDB
	//outputs: 2 outputs; 1 is reg number, 1 is data
);

//Process to reorder

endmodule